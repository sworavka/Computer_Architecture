module singlecycle(
    input resetl,
    input [63:0] startpc,
    output reg [63:0] currentpc,
    output [63:0] dmemout,
    input CLK
);

    // Next PC connections
    wire [63:0] nextpc;       // The next PC, to be updated on clock cycle

    // Instruction Memory connections
    wire [31:0] instruction;  // The current instruction

    // Parts of instruction
    wire [4:0] rd;            // The destination register
    wire [4:0] rm;            // Operand 1
    wire [4:0] rn;            // Operand 2
    wire [10:0] opcode;

    // Control wires
    wire reg2loc;
    wire alusrc;
    wire mem2reg;
    wire regwrite;
    wire memread;
    wire memwrite;
    wire branch;
    wire uncond_branch;
    wire [3:0] aluctrl;
    wire [1:0] signop;

    // Register file connections
    wire [63:0] regoutA;     // Output A
    wire [63:0] regoutB;     // Output B

    // ALU connections
    wire [63:0] aluout;
    wire zero;

    // Sign Extender connections
    wire [63:0] extimm;

    // PC update logic
    always @(negedge CLK)
    begin
        if (resetl)
            currentpc <= nextpc;
        else
            currentpc <= startpc;
    end

    // Parts of instruction
    assign rd = instruction[4:0];
    assign rm = instruction[9:5];
    assign rn = reg2loc ? instruction[4:0] : instruction[20:16];
    assign opcode = instruction[31:21];

    // Instruction Memory
    InstructionMemory imem(
        .Data(instruction),
        .Address(currentpc)
    );

    // Control Unit
    control control(
        .reg2loc(reg2loc),
        .alusrc(alusrc),
        .mem2reg(mem2reg),
        .regwrite(regwrite),
        .memread(memread),
        .memwrite(memwrite),
        .branch(branch),
        .uncond_branch(uncond_branch),
        .aluop(aluctrl),
        .signop(signop),
        .opcode(opcode)
    );

    // Register File
    RegisterFile regfile(
        .ReadReg1(rn),
        .ReadReg2(rm),
        .WriteReg(rd),
        .WriteData(dmemout),
        .RegWrite(regwrite),
        .ReadData1(regoutA),
        .ReadData2(regoutB),
        .Clk(CLK)
    );

    // ALU
    ALU alu(
        .ALUControl(aluctrl),
        .A(regoutA),
        .B(alusrc ? extimm : regoutB),
        .ALUResult(aluout),
        .Zero(zero)
    );

    // Sign Extender
    SignExtender signext(
        .SignOp(signop),
        .Instr(instruction[20:0]),
        .Out(extimm)
    );

    // Data Memory
    DataMemory dmem(
        .Address(aluout),
        .WriteData(regoutB),
        .ReadData(dmemout),
        .MemWrite(memwrite),
        .MemRead(memread),
        .Clk(CLK)
    );

    // Next PC logic
    assign nextpc = (uncond_branch || (branch && zero)) ? (currentpc + (extimm << 2)) : (currentpc + 4);

endmodule
